/////////////////////////////////////////////
// aes
//   Top level module with SPI interface and SPI core
/////////////////////////////////////////////

module aes_cipher(input  logic clk,
           input  logic sck, 
           input  logic sdi,
           output logic sdo,
           input  logic load,
           output logic done);
                    
    logic [127:0] key, plaintext, cyphertext;
            
    aes_spi spi(sck, sdi, sdo, done, key, plaintext, cyphertext);   
    aes_core core(clk, load, key, plaintext, done, cyphertext);
endmodule

/////////////////////////////////////////////
// aes_spi
//   SPI interface.  Shifts in key and plaintext
//   Captures ciphertext when done, then shifts it out
//   Tricky cases to properly change sdo on negedge clk
/////////////////////////////////////////////

module aes_spi(input  logic sck, 
               input  logic sdi,
               output logic sdo,
               input  logic done,
               output logic [127:0] key, plaintext,
               input  logic [127:0] cyphertext);

    logic         sdodelayed, wasdone;
    logic [127:0] cyphertextcaptured;
               
    // assert load
    // apply 256 sclks to shift in key and plaintext, starting with plaintext[127]
    // then deassert load, wait until done
    // then apply 128 sclks to shift out cyphertext, starting with cyphertext[127]
    // SPI mode is equivalent to cpol = 0, cpha = 0 since data is sampled on first edge and the first
    // edge is a rising edge (clock going from low in the idle state to high).
    always_ff @(posedge sck)
        if (!wasdone)  {cyphertextcaptured, plaintext, key} = {cyphertext, plaintext[126:0], key, sdi};
        else           {cyphertextcaptured, plaintext, key} = {cyphertextcaptured[126:0], plaintext, key, sdi}; 
    
    // sdo should change on the negative edge of sck
    always_ff @(negedge sck) begin
        wasdone = done;
        sdodelayed = cyphertextcaptured[126];
    end
    
    // when done is first asserted, shift out msb before clock edge
    assign sdo = (done & !wasdone) ? cyphertext[127] : sdodelayed;
endmodule

/////////////////////////////////////////////
// aes_core
//   top level AES encryption module
//   when load is asserted, takes the current key and plaintext
//   generates cyphertext and asserts done when complete 11 cycles later
// 
//   See FIPS-197 with Nk = 4, Nb = 4, Nr = 10
//
//   The key and message are 128-bit values packed into an array of 16 bytes as
//   shown below
//        [127:120] [95:88] [63:56] [31:24]     S0,0    S0,1    S0,2    S0,3
//        [119:112] [87:80] [55:48] [23:16]     S1,0    S1,1    S1,2    S1,3
//        [111:104] [79:72] [47:40] [15:8]      S2,0    S2,1    S2,2    S2,3
//        [103:96]  [71:64] [39:32] [7:0]       S3,0    S3,1    S3,2    S3,3
//
//   Equivalently, the values are packed into four words as given
//        [127:96]  [95:64] [63:32] [31:0]      w[0]    w[1]    w[2]    w[3]
/////////////////////////////////////////////

module aes_core(input  logic         clk,
                input  logic         load,
                input  logic [127:0] key, 
                input  logic [127:0] plaintext, 
                output logic         done, 
                output logic [127:0] cyphertext);
    // TODO: Your code goes here
	logic [127:0] firststate, prevstate, state;
	logic counter;
	logic [3:0] round;

	always_ff @(posedge clk) begin
		if (load == 0) begin
			counter <= 1'b0;
			round <= 4'b0;
		end
		else if (counter[1] == 1) begin
			counter <= counter + 1;
			round <= round + 1;
		end
		else		begin
			counter <= counter + 1;
			round <= round;
		end
	end

	assign mux1 = ((round==4'd0) | (round == 4'd9)) ? state_after_firstaddkey : state_after_addkey;
	assign mux2 = (round == 4'd9) ? state : prevstate;
	assign prevstate = mux2;

	addroundkey(state, key, state_after_firstaddkey);
	findnextkey(key, round, nextkey);
	subbytes(mux1, state_after_subbytes);
	shiftrows(state_after_subbytes, state_after_shiftrows);
	mixcolumns(state_after_shiftrows, state_after_mixcols);
	addroundkey(state_after_mixcols, nextkey, state_after_addkey);

	findnextkey(key, round, key)
	subbytes(mux2, state);
	shiftrows(state, state);
	addroundkey(state, key, state);

	assign cyphertext = state;
	
	
    
endmodule

/////////////////////////////////////////////
// addroundkey
//   Infamous AES byte substitutions with magic numbers
//   Combinational version which is mapped to LUTs (logic cells)
//   Section 5.1.4
/////////////////////////////////////////////
module addroundkey(input logic [127:0] a,
				   input logic [127:0] key,
				   output logic [127:0] y);
	assign y = a ^ key; 
endmodule

/////////////////////////////////////////////
// findnextkey
//   Figures out what the next key is based on current round and current key
//   The next key is the next column of the input keys
/////////////////////////////////////////////
module findnextkey(input logic [127:0] prevkey,
				   input logic [3:0] round,
				   output logic [127:0] nextkey);
	logic [31:0] rcon;
	logic [31:0] rotword;
	logic [7:0] subbytes1, subbytes2, subbytes3, subbytes4;
	logic [31:0] subbytes;
	logic [31:0] firstcol seccol, thirdcol, fourcol;
	assign rotword = {prevkey[23:0], prevkey[31:24]};
	
	sbox_sync(rotword[31:24], subbytes1);
	sbox_sync(rotword[23:16], subbytes2);
	sbox_sync(rotword[15:8], subbytes3);
	sbox_sync(rotword[7:0], subbytes4);

	assign subbytes = {subbytes1, subbytes2, subbytes3, subbytes4};
	
	always_comb begin
		case (round)
			4'd1:		rcon = {8'h01, 24'h0};
			4'd2:		rcon = {8'h02, 24'h0};
			4'd3:		rcon = {8'h04, 24'h0};
			4'd4:		rcon = {8'h08, 24'h0};
			4'd5:		rcon = {8'h10, 24'h0};
			4'd6:		rcon = {8'h20, 24'h0};
			4'd7:		rcon = {8'h40, 24'h0};
			4'd8:		rcon = {8'h80, 24'h0};
			4'd9:		rcon = {8'h1b, 24'h0};
			4'd10:		rcon = {8'h36, 24'h0};
			default: 	rcon = 32'h0;
		endcase
	end	

	assign firstcol = key[127:96] ^ subbytes ^ rotword;
	assign seccol = key[95:64] ^ firstcol;
	assign thirdcol = key[63:32] ^ seccol;
	assign fourcol = key[31:0] ^ thirdcol;
	assign nextkey = {firstcol, seccol, thirdcol, fourcol};
endmodule

/////////////////////////////////////////////
// sbox
//   Infamous AES byte substitutions with magic numbers
//   Combinational version which is mapped to LUTs (logic cells)
//   Section 5.1.1, Figure 7
/////////////////////////////////////////////

module sbox(input  logic [7:0] a,
            output logic [7:0] y);
            
  // sbox implemented as a ROM
  // This module is combinational and will be inferred using LUTs (logic cells)
  logic [7:0] sbox[0:255];

  initial   $readmemh("sbox.txt", sbox);
  assign y = sbox[a];
endmodule

/////////////////////////////////////////////
// subbytes
//   AES byte substitution for the whole text
//   Uses synchronous sbox
//   Section 5.1.1
/////////////////////////////////////////////
module subbytes(
	input		logic [127:0] a,
	output 	logic [127:0] y);
            
  // sbox implemented as a ROM
  // This module is synchronous and will be inferred using BRAMs (Block RAMs)
	sbox_sync(a[127:120], y[127:120]);
	sbox_sync(a[119:112], y[119:112]);
	sbox_sync(a[111:104], y[111:104]);
	sbox_sync(a[103:96], y[103:96]);
	sbox_sync(a[95:88], y[95:88]);
	sbox_sync(a[87:80], y[87:80]);
	sbox_sync(a[79:72], y[79:72]);
	sbox_sync(a[71:64], y[71:64]);
	sbox_sync(a[63:56], y[63:56]);
	sbox_sync(a[55:48], y[55:48]);
	sbox_sync(a[47:40], y[47:40]);
	sbox_sync(a[39:32], y[39:32]);
	sbox_sync(a[31:24], y[31:24]);
	sbox_sync(a[23:16], y[23:16]);
	sbox_sync(a[15:8], y[15:8]);
	sbox_sync(a[7:0], y[7:0]);
endmodule

/////////////////////////////////////////////
// sbox
//   Infamous AES byte substitutions with magic numbers
//   Synchronous version which is mapped to embedded block RAMs (EBR)
//   Section 5.1.1, Figure 7
/////////////////////////////////////////////
module sbox_sync(
	input		logic [7:0] a,
	input	 	logic 			clk,
	output 	logic [7:0] y);
            
  // sbox implemented as a ROM
  // This module is synchronous and will be inferred using BRAMs (Block RAMs)
  logic [7:0] sbox [0:255];

  initial   $readmemh("sbox.txt", sbox);
	
	// Synchronous version
	always_ff @(posedge clk) begin
		y <= sbox[a];
	end
endmodule

/////////////////////////////////////////////
// shiftrows
//   The bytes in the last three rows of the State are cyclically shifted over different numbers of bytes
//   Section 5.1.2, Figure 8
//   Operation different for each row, use array swizzling
/////////////////////////////////////////////

module shiftrows(input  logic [127:0] a,
                 output logic [127:0] y);
	assign y = {a[127:120], a[87:80], a[47:40], a[7:0],
				a[95:88], a[55:48], a[15:8], a[103:96],
				a[63:56], a[23:16], a[111:104], a[71:64],
				a[31:24], a[119:112], a[79:72], a[39:32]}
endmodule

/////////////////////////////////////////////
// mixcolumns
//   Even funkier action on columns
//   Section 5.1.3, Figure 9
//   Same operation performed on each of four columns
/////////////////////////////////////////////

module mixcolumns(input  logic [127:0] a,
                  output logic [127:0] y);

  mixcolumn mc0(a[127:96], y[127:96]);
  mixcolumn mc1(a[95:64],  y[95:64]);
  mixcolumn mc2(a[63:32],  y[63:32]);
  mixcolumn mc3(a[31:0],   y[31:0]);
endmodule

/////////////////////////////////////////////
// mixcolumn
//   Perform Galois field operations on bytes in a column
//   See EQ(4) from E. Ahmed et al, Lightweight Mix Columns Implementation for AES, AIC09
//   for this hardware implementation
/////////////////////////////////////////////

module mixcolumn(input  logic [31:0] a,
                 output logic [31:0] y);
                      
        logic [7:0] a0, a1, a2, a3, y0, y1, y2, y3, t0, t1, t2, t3, tmp;
        
        assign {a0, a1, a2, a3} = a;
        assign tmp = a0 ^ a1 ^ a2 ^ a3;
    
        galoismult gm0(a0^a1, t0);
        galoismult gm1(a1^a2, t1);
        galoismult gm2(a2^a3, t2);
        galoismult gm3(a3^a0, t3);
        
        assign y0 = a0 ^ tmp ^ t0;
        assign y1 = a1 ^ tmp ^ t1;
        assign y2 = a2 ^ tmp ^ t2;
        assign y3 = a3 ^ tmp ^ t3;
        assign y = {y0, y1, y2, y3};    
endmodule

/////////////////////////////////////////////
// galoismult
//   Multiply by x in GF(2^8) is a left shift
//   followed by an XOR if the result overflows
//   Uses irreducible polynomial x^8+x^4+x^3+x+1 = 00011011
/////////////////////////////////////////////

module galoismult(input  logic [7:0] a,
                  output logic [7:0] y);

    logic [7:0] ashift;
    
    assign ashift = {a[6:0], 1'b0};
    assign y = a[7] ? (ashift ^ 8'b00011011) : ashift;
endmodule
